library verilog;
use verilog.vl_types.all;
entity SimpleCompArch_vlg_vec_tst is
end SimpleCompArch_vlg_vec_tst;
